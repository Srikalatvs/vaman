module sevenseg(output a, output b,output c,output d,output e,output f,output g);
assign a = 0;
assign b = 0;
assign c = 0;
assign d = 0;
assign e = 0;
assign f = 0;
assign g = 1;
endmodule
   
